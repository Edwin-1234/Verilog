module nor_gate(input a,b,output y);
  nor(y,a,b);
endmodule
