module not_gate(input x,output y);
  not(y,x);
endmodule
